/*
 * =====================================================================
 * (c) Copyright 2001  BBNT Solutions, LLC
 * =====================================================================
 */

contract Logging ( )
{
    region Normal (true ) 
	{}
};

