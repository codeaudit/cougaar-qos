/*
 * =====================================================================
 * (c) Copyright 2001  BBNT Solutions, LLC
 * =====================================================================
 */

contract RemoteSSL
    (
     syscond quo::ExpectedCapacitySC quo_data::ExpectedCapacitySCImpl Bandwidth,
     syscond quo::ValueSC ValueSCImpl UseSSL,

     syscond quo::ValueSC ValueSCImpl trust
     
     )
{
  region ForceSSL (UseSSL )
    {}
  region AdaptiveSSL (true) {
    region Compromised (trust == 0) {
      region SameHost (Bandwidth >= 1000000)
	{}
      region SameLan  (Bandwidth >= 10000)
	{}
      region Wan  (true)  
	{}
    }
    region Suspect (trust <= 2) {
      region SameHost (Bandwidth >= 10000000)
	{}
      region SameLan  (Bandwidth >= 10000)
	{}
      region Wan  (true)  
	{}
    }
    region Normal (trust <= 5) {
      region SameHost (Bandwidth >= 10000000)
	{}
      region SameLan  (Bandwidth >= 10000)
	{}
      region Wan  (true)  
	{}
    }
    region CareFree (trust <= 10) {
      region SameHost (Bandwidth >= 10000000)
	{}
      region SameLan  (Bandwidth >= 10000)
	{}
      region Wan  (true)  
	{}
    }
  }
};
