/*
 * =====================================================================
 * (c) Copyright 2001  BBNT Solutions, LLC
 * =====================================================================
 */

contract Diagnose  ()
{
  region Normal (true) {}

};

